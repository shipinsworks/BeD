`ifndef _C2SIF_SVH_
 `define _C2SIF_SVH_

 `include "macro.svh"

interface c2sif();
   
endinterface // c2sif

`endif
