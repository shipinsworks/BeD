`ifndef _DPI_C_SVH_
 `define _DPI_C_SVH_

   import "DPI-C" context task scenario();
   export "DPI-C" task cs_printf;
   
`endif
