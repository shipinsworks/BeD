`ifndef _MACRO_SVH_
 `define _MACRO_SVH_

 `define debug_printf( msg ) $display( "[Debug   ] %8d : %s", $stime, $sformatf( msg ))

`endif
